library verilog;
use verilog.vl_types.all;
entity bcdAdd_vlg_vec_tst is
end bcdAdd_vlg_vec_tst;
