library verilog;
use verilog.vl_types.all;
entity \1fa\ is
    port(
        S               : out    vl_logic;
        Ci              : in     vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        Co              : out    vl_logic
    );
end \1fa\;
